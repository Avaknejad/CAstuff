library verilog;
use verilog.vl_types.all;
entity MultiplierTest is
end MultiplierTest;
